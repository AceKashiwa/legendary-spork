`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/19 13:42:37
// Design Name: 
// Module Name: ssd1306_spi4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ssd1306_spi4(
    input clk,
    input rst_n,
    output oled_rst_n,  // RES
    output oled_cs_n,   // CS
    output oled_dc,     // DC
    output oled_clk,    // SCL  D0
    output oled_data    // SDA  D1
    );
    

endmodule
