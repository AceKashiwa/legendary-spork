`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/24
// Design Name: 
// Module Name: music_score_ROM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 乐谱信息ROM，每一节拍输出音符编码，只读优化版
// 
//////////////////////////////////////////////////////////////////////////////////

module music_score_ROM #(
    parameter ROM_WIDTH = 12,      // {high[3:0], med[3:0], low[3:0]}
    parameter ROM_DEPTH = 135,     // 节拍数
    parameter ADDR_WIDTH = 8
)(
    input [ADDR_WIDTH-1:0] addr,
    output reg [ROM_WIDTH-1:0] data
);
    reg [ROM_WIDTH-1:0] Mem[ROM_DEPTH-1:0];

    // 初始化ROM内容
    initial begin
        // {high, med, low}
        Mem[  0] = {4'h0, 4'h0, 4'h3};
        Mem[  1] = {4'h0, 4'h0, 4'h3};
        Mem[  2] = {4'h0, 4'h0, 4'h3};
        Mem[  3] = {4'h0, 4'h0, 4'h3};
        Mem[  4] = {4'h0, 4'h0, 4'h5};
        Mem[  5] = {4'h0, 4'h0, 4'h5};
        Mem[  6] = {4'h0, 4'h0, 4'h5};
        Mem[  7] = {4'h0, 4'h0, 4'h6};
        Mem[  8] = {4'h0, 4'h1, 4'h0};
        Mem[  9] = {4'h0, 4'h1, 4'h0};
        Mem[ 10] = {4'h0, 4'h1, 4'h0};
        Mem[ 11] = {4'h0, 4'h2, 4'h0};
        Mem[ 12] = {4'h0, 4'h0, 4'h6};
        Mem[ 13] = {4'h0, 4'h1, 4'h0};
        Mem[ 14] = {4'h0, 4'h0, 4'h5};
        Mem[ 15] = {4'h0, 4'h0, 4'h5};

        Mem[ 16] = {4'h0, 4'h5, 4'h0};
        Mem[ 17] = {4'h0, 4'h5, 4'h0};
        Mem[ 18] = {4'h0, 4'h5, 4'h0};
        Mem[ 19] = {4'h1, 4'h0, 4'h0};
        Mem[ 20] = {4'h0, 4'h6, 4'h0};
        Mem[ 21] = {4'h0, 4'h5, 4'h0};
        Mem[ 22] = {4'h0, 4'h3, 4'h0};
        Mem[ 23] = {4'h0, 4'h5, 4'h0};
        Mem[ 24] = {4'h0, 4'h2, 4'h0};
        Mem[ 25] = {4'h0, 4'h2, 4'h0};
        Mem[ 26] = {4'h0, 4'h2, 4'h0};
        Mem[ 27] = {4'h0, 4'h2, 4'h0};
        Mem[ 28] = {4'h0, 4'h2, 4'h0};
        Mem[ 29] = {4'h0, 4'h2, 4'h0};
        Mem[ 30] = {4'h0, 4'h0, 4'h0};
        Mem[ 31] = {4'h0, 4'h0, 4'h0};

        Mem[ 32] = {4'h0, 4'h2, 4'h0};
        Mem[ 33] = {4'h0, 4'h2, 4'h0};
        Mem[ 34] = {4'h0, 4'h2, 4'h0};
        Mem[ 35] = {4'h0, 4'h3, 4'h0};
        Mem[ 36] = {4'h0, 4'h0, 4'h7};
        Mem[ 37] = {4'h0, 4'h0, 4'h7};
        Mem[ 38] = {4'h0, 4'h0, 4'h6};
        Mem[ 39] = {4'h0, 4'h0, 4'h6};
        Mem[ 40] = {4'h0, 4'h0, 4'h5};
        Mem[ 41] = {4'h0, 4'h0, 4'h5};
        Mem[ 42] = {4'h0, 4'h0, 4'h5};
        Mem[ 43] = {4'h0, 4'h0, 4'h6};
        Mem[ 44] = {4'h0, 4'h1, 4'h0};
        Mem[ 45] = {4'h0, 4'h1, 4'h0};
        Mem[ 46] = {4'h0, 4'h2, 4'h0};
        Mem[ 47] = {4'h0, 4'h2, 4'h0};

        Mem[ 48] = {4'h0, 4'h0, 4'h3};
        Mem[ 49] = {4'h0, 4'h0, 4'h3};
        Mem[ 50] = {4'h0, 4'h1, 4'h0};
        Mem[ 51] = {4'h0, 4'h1, 4'h0};
        Mem[ 52] = {4'h0, 4'h0, 4'h6};
        Mem[ 53] = {4'h0, 4'h0, 4'h5};
        Mem[ 54] = {4'h0, 4'h0, 4'h6};
        Mem[ 55] = {4'h0, 4'h1, 4'h0};
        Mem[ 56] = {4'h0, 4'h0, 4'h5};
        Mem[ 57] = {4'h0, 4'h0, 4'h5};
        Mem[ 58] = {4'h0, 4'h0, 4'h5};
        Mem[ 59] = {4'h0, 4'h0, 4'h5};
        Mem[ 60] = {4'h0, 4'h0, 4'h5};
        Mem[ 61] = {4'h0, 4'h0, 4'h5};
        Mem[ 62] = {4'h0, 4'h0, 4'h5};
        Mem[ 63] = {4'h0, 4'h0, 4'h5};

        Mem[ 64] = {4'h0, 4'h3, 4'h0};
        Mem[ 65] = {4'h0, 4'h3, 4'h0};
        Mem[ 66] = {4'h0, 4'h3, 4'h0};
        Mem[ 67] = {4'h0, 4'h5, 4'h0};
        Mem[ 68] = {4'h0, 4'h0, 4'h7};
        Mem[ 69] = {4'h0, 4'h0, 4'h7};
        Mem[ 70] = {4'h0, 4'h2, 4'h0};
        Mem[ 71] = {4'h0, 4'h2, 4'h0};
        Mem[ 72] = {4'h0, 4'h0, 4'h6};
        Mem[ 73] = {4'h0, 4'h1, 4'h0};
        Mem[ 74] = {4'h0, 4'h0, 4'h5};
        Mem[ 75] = {4'h0, 4'h0, 4'h5};
        Mem[ 76] = {4'h0, 4'h0, 4'h5};
        Mem[ 77] = {4'h0, 4'h0, 4'h5};
        Mem[ 78] = {4'h0, 4'h0, 4'h0};
        Mem[ 79] = {4'h0, 4'h0, 4'h0};

        Mem[ 80] = {4'h0, 4'h0, 4'h3};
        Mem[ 81] = {4'h0, 4'h0, 4'h5};
        Mem[ 82] = {4'h0, 4'h0, 4'h5};
        Mem[ 83] = {4'h0, 4'h0, 4'h3};
        Mem[ 84] = {4'h0, 4'h0, 4'h5};
        Mem[ 85] = {4'h0, 4'h0, 4'h6};
        Mem[ 86] = {4'h0, 4'h0, 4'h7};
        Mem[ 87] = {4'h0, 4'h2, 4'h0};
        Mem[ 88] = {4'h0, 4'h0, 4'h6};
        Mem[ 89] = {4'h0, 4'h0, 4'h6};
        Mem[ 90] = {4'h0, 4'h0, 4'h6};
        Mem[ 91] = {4'h0, 4'h0, 4'h6};
        Mem[ 92] = {4'h0, 4'h0, 4'h6};
        Mem[ 93] = {4'h0, 4'h0, 4'h6};
        Mem[ 94] = {4'h0, 4'h0, 4'h5};
        Mem[ 95] = {4'h0, 4'h0, 4'h6};

        Mem[ 96] = {4'h0, 4'h1, 4'h0};
        Mem[ 97] = {4'h0, 4'h1, 4'h0};
        Mem[ 98] = {4'h0, 4'h1, 4'h0};
        Mem[ 99] = {4'h0, 4'h2, 4'h0};
        Mem[100] = {4'h0, 4'h5, 4'h0};
        Mem[101] = {4'h0, 4'h5, 4'h0};
        Mem[102] = {4'h0, 4'h3, 4'h0};
        Mem[103] = {4'h0, 4'h3, 4'h0};
        Mem[104] = {4'h0, 4'h2, 4'h0};
        Mem[105] = {4'h0, 4'h2, 4'h0};
        Mem[106] = {4'h0, 4'h3, 4'h0};
        Mem[107] = {4'h0, 4'h2, 4'h0};
        Mem[108] = {4'h0, 4'h1, 4'h0};
        Mem[109] = {4'h0, 4'h1, 4'h0};
        Mem[110] = {4'h0, 4'h0, 4'h6};
        Mem[111] = {4'h0, 4'h0, 4'h5};

        Mem[112] = {4'h0, 4'h0, 4'h3};
        Mem[113] = {4'h0, 4'h0, 4'h3};
        Mem[114] = {4'h0, 4'h0, 4'h3};
        Mem[115] = {4'h0, 4'h0, 4'h3};
        Mem[116] = {4'h0, 4'h1, 4'h0};
        Mem[117] = {4'h0, 4'h1, 4'h0};
        Mem[118] = {4'h0, 4'h1, 4'h0};
        Mem[119] = {4'h0, 4'h1, 4'h0};
        Mem[120] = {4'h0, 4'h0, 4'h6};
        Mem[121] = {4'h0, 4'h1, 4'h0};
        Mem[122] = {4'h0, 4'h0, 4'h6};
        Mem[123] = {4'h0, 4'h0, 4'h5};
        Mem[124] = {4'h0, 4'h0, 4'h3};
        Mem[125] = {4'h0, 4'h0, 4'h5};
        Mem[126] = {4'h0, 4'h0, 4'h6};
        Mem[127] = {4'h0, 4'h1, 4'h0};

        Mem[128] = {4'h0, 4'h0, 4'h5};
        Mem[129] = {4'h0, 4'h0, 4'h5};
        Mem[130] = {4'h0, 4'h0, 4'h5};
        Mem[131] = {4'h0, 4'h0, 4'h5};
        Mem[132] = {4'h0, 4'h0, 4'h5};
        Mem[133] = {4'h0, 4'h0, 4'h0};
        Mem[134] = {4'h0, 4'h0, 4'h0};
    end

    always @(*) begin
        data = Mem[addr];
    end

endmodule