`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/24
// Design Name: 
// Module Name: music_score_ROM_xxx
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 小星星乐谱ROM，只读、组合逻辑输出
// 
//////////////////////////////////////////////////////////////////////////////////

module music_score_ROM_xxx #(
    parameter ROM_WIDTH = 12,      // {high[3:0], med[3:0], low[3:0]}
    parameter ROM_DEPTH = 96,    // 96音符
    parameter ADDR_WIDTH = 7
)(
    input  [ADDR_WIDTH-1:0] addr,
    output [ROM_WIDTH-1:0]  data
);
    reg [ROM_WIDTH-1:0] Mem[0:ROM_DEPTH-1];

    // 小星星简谱：1 1 5 5 6 6 5 | 4 4 3 3 2 2 1 | 5 5 4 4 3 3 2 | 5 5 4 4 3 3 2 | 1 1 5 5 6 6 5 | 4 4 3 3 2 2 1
    // 只用C调，1=C，2=D，3=E，4=F，5=G，6=A
    // 低音：{4'h0, 4'h0, 4'hX}，X为音符
    // 静音：{4'h0, 4'h0, 4'h0}
    initial begin
        Mem[ 0] = {4'h0, 4'h0, 4'h1}; // 1
        Mem[ 1] = {4'h0, 4'h0, 4'h1}; // 1
        Mem[ 2] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[ 3] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[ 4] = {4'h0, 4'h0, 4'h6}; // 6
        Mem[ 5] = {4'h0, 4'h0, 4'h6}; // 6
        Mem[ 6] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[ 7] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[ 8] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[ 9] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[10] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[11] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[12] = {4'h0, 4'h0, 4'h2}; // 2
        Mem[13] = {4'h0, 4'h0, 4'h2}; // 2
        Mem[14] = {4'h0, 4'h0, 4'h1}; // 1
        Mem[15] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[16] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[17] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[18] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[19] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[20] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[21] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[22] = {4'h0, 4'h0, 4'h2}; // 2
        Mem[23] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[24] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[25] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[26] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[27] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[28] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[29] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[30] = {4'h0, 4'h0, 4'h2}; // 2
        Mem[31] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[32] = {4'h0, 4'h0, 4'h1}; // 1
        Mem[33] = {4'h0, 4'h0, 4'h1}; // 1
        Mem[34] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[35] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[36] = {4'h0, 4'h0, 4'h6}; // 6
        Mem[37] = {4'h0, 4'h0, 4'h6}; // 6
        Mem[38] = {4'h0, 4'h0, 4'h5}; // 5
        Mem[39] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[40] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[41] = {4'h0, 4'h0, 4'h4}; // 4
        Mem[42] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[43] = {4'h0, 4'h0, 4'h3}; // 3
        Mem[44] = {4'h0, 4'h0, 4'h2}; // 2
        Mem[45] = {4'h0, 4'h0, 4'h2}; // 2
        Mem[46] = {4'h0, 4'h0, 4'h1}; // 1
        Mem[47] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）
        // 升调
        Mem[48] = {4'h0, 4'h1, 4'h0}; // 1
        Mem[49] = {4'h0, 4'h1, 4'h0}; // 1
        Mem[50] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[51] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[52] = {4'h0, 4'h6, 4'h0}; // 6
        Mem[53] = {4'h0, 4'h6, 4'h0}; // 6
        Mem[54] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[55] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[56] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[57] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[58] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[59] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[60] = {4'h0, 4'h2, 4'h0}; // 2
        Mem[61] = {4'h0, 4'h2, 4'h0}; // 2
        Mem[62] = {4'h0, 4'h1, 4'h0}; // 1
        Mem[63] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[64] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[65] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[66] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[67] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[68] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[69] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[70] = {4'h0, 4'h2, 4'h0}; // 2
        Mem[71] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[72] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[73] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[74] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[75] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[76] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[77] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[78] = {4'h0, 4'h2, 4'h0}; // 2
        Mem[79] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[80] = {4'h0, 4'h1, 4'h0}; // 1
        Mem[81] = {4'h0, 4'h1, 4'h0}; // 1
        Mem[82] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[83] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[84] = {4'h0, 4'h6, 4'h0}; // 6
        Mem[85] = {4'h0, 4'h6, 4'h0}; // 6
        Mem[86] = {4'h0, 4'h5, 4'h0}; // 5
        Mem[87] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）

        Mem[88] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[89] = {4'h0, 4'h4, 4'h0}; // 4
        Mem[90] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[91] = {4'h0, 4'h3, 4'h0}; // 3
        Mem[92] = {4'h0, 4'h2, 4'h0}; // 2
        Mem[93] = {4'h0, 4'h2, 4'h0}; // 2
        Mem[94] = {4'h0, 4'h1, 4'h0}; // 1
        Mem[95] = {4'h0, 4'h0, 4'h0}; // |（间隔或延音）
        end

    assign data = Mem[addr];

endmodule