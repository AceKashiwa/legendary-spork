`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/24
// Design Name: 
// Module Name: music_score_ROM_xxx
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 小星星乐谱ROM
// 
//////////////////////////////////////////////////////////////////////////////////

module music_score_ROM_xxx #(
    parameter ROM_WIDTH = 12,      // {high[3:0], med[3:0], low[3:0]}
    parameter ROM_DEPTH = 128,     // 128拍
    parameter ADDR_WIDTH = 7
)(
    input  [ADDR_WIDTH-1:0] addr,
    output [ROM_WIDTH-1:0]  data
);
    reg [ROM_WIDTH-1:0] Mem[0:ROM_DEPTH-1];

    // 1 1 5 5 6 6 5 0
    // 4 4 3 3 2 2 1 0
    // 5 5 4 4 3 3 2 0
    // 5 5 4 4 3 3 2 0
    initial begin
        Mem[  0] = {4'h0, 4'h0, 4'h1};
        Mem[  1] = {4'h0, 4'h0, 4'h1};
        Mem[  2] = {4'h0, 4'h0, 4'h1};
        Mem[  3] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[  4] = {4'h0, 4'h0, 4'h1};
        Mem[  5] = {4'h0, 4'h0, 4'h1};
        Mem[  6] = {4'h0, 4'h0, 4'h1};
        Mem[  7] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[  8] = {4'h0, 4'h0, 4'h5};
        Mem[  9] = {4'h0, 4'h0, 4'h5};
        Mem[ 10] = {4'h0, 4'h0, 4'h5};
        Mem[ 11] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 12] = {4'h0, 4'h0, 4'h5};
        Mem[ 13] = {4'h0, 4'h0, 4'h5};
        Mem[ 14] = {4'h0, 4'h0, 4'h5};
        Mem[ 15] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 16] = {4'h0, 4'h0, 4'h6};
        Mem[ 17] = {4'h0, 4'h0, 4'h6};
        Mem[ 18] = {4'h0, 4'h0, 4'h6};
        Mem[ 19] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 20] = {4'h0, 4'h0, 4'h6};
        Mem[ 21] = {4'h0, 4'h0, 4'h6};
        Mem[ 22] = {4'h0, 4'h0, 4'h6};
        Mem[ 23] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 24] = {4'h0, 4'h0, 4'h5};
        Mem[ 25] = {4'h0, 4'h0, 4'h5};
        Mem[ 26] = {4'h0, 4'h0, 4'h5};
        Mem[ 27] = {4'h0, 4'h0, 4'h5};
        Mem[ 28] = {4'h0, 4'h0, 4'h5};
        Mem[ 29] = {4'h0, 4'h0, 4'h5};
        Mem[ 30] = {4'h0, 4'h0, 4'h5};
        Mem[ 31] = {4'h0, 4'h0, 4'h0}; // 空

        Mem[ 32] = {4'h0, 4'h0, 4'h4};
        Mem[ 33] = {4'h0, 4'h0, 4'h4};
        Mem[ 34] = {4'h0, 4'h0, 4'h4};
        Mem[ 35] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 36] = {4'h0, 4'h0, 4'h4};
        Mem[ 37] = {4'h0, 4'h0, 4'h4};
        Mem[ 38] = {4'h0, 4'h0, 4'h4};
        Mem[ 39] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 40] = {4'h0, 4'h0, 4'h3};
        Mem[ 41] = {4'h0, 4'h0, 4'h3};
        Mem[ 42] = {4'h0, 4'h0, 4'h3};
        Mem[ 43] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 44] = {4'h0, 4'h0, 4'h3};
        Mem[ 45] = {4'h0, 4'h0, 4'h3};
        Mem[ 46] = {4'h0, 4'h0, 4'h3};
        Mem[ 47] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 48] = {4'h0, 4'h0, 4'h2};
        Mem[ 49] = {4'h0, 4'h0, 4'h2};
        Mem[ 50] = {4'h0, 4'h0, 4'h2};
        Mem[ 51] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 52] = {4'h0, 4'h0, 4'h2};
        Mem[ 53] = {4'h0, 4'h0, 4'h2};
        Mem[ 54] = {4'h0, 4'h0, 4'h2};
        Mem[ 55] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 56] = {4'h0, 4'h0, 4'h1};
        Mem[ 57] = {4'h0, 4'h0, 4'h1};
        Mem[ 58] = {4'h0, 4'h0, 4'h1};
        Mem[ 59] = {4'h0, 4'h0, 4'h1};
        Mem[ 60] = {4'h0, 4'h0, 4'h1};
        Mem[ 61] = {4'h0, 4'h0, 4'h1};
        Mem[ 62] = {4'h0, 4'h0, 4'h1};
        Mem[ 63] = {4'h0, 4'h0, 4'h0}; // 空

        Mem[ 64] = {4'h0, 4'h0, 4'h5};
        Mem[ 65] = {4'h0, 4'h0, 4'h5};
        Mem[ 66] = {4'h0, 4'h0, 4'h5};
        Mem[ 67] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 68] = {4'h0, 4'h0, 4'h5};
        Mem[ 69] = {4'h0, 4'h0, 4'h5};
        Mem[ 70] = {4'h0, 4'h0, 4'h5};
        Mem[ 71] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 72] = {4'h0, 4'h0, 4'h4};
        Mem[ 73] = {4'h0, 4'h0, 4'h4};
        Mem[ 74] = {4'h0, 4'h0, 4'h4};
        Mem[ 75] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 76] = {4'h0, 4'h0, 4'h4};
        Mem[ 77] = {4'h0, 4'h0, 4'h4};
        Mem[ 78] = {4'h0, 4'h0, 4'h4};
        Mem[ 79] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 80] = {4'h0, 4'h0, 4'h3};
        Mem[ 81] = {4'h0, 4'h0, 4'h3};
        Mem[ 82] = {4'h0, 4'h0, 4'h3};
        Mem[ 83] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 84] = {4'h0, 4'h0, 4'h3};
        Mem[ 85] = {4'h0, 4'h0, 4'h3};
        Mem[ 86] = {4'h0, 4'h0, 4'h3};
        Mem[ 87] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[ 88] = {4'h0, 4'h0, 4'h2};
        Mem[ 89] = {4'h0, 4'h0, 4'h2};
        Mem[ 90] = {4'h0, 4'h0, 4'h2};
        Mem[ 91] = {4'h0, 4'h0, 4'h2};
        Mem[ 92] = {4'h0, 4'h0, 4'h2};
        Mem[ 93] = {4'h0, 4'h0, 4'h2};
        Mem[ 94] = {4'h0, 4'h0, 4'h2};
        Mem[ 95] = {4'h0, 4'h0, 4'h0}; // 空
        
        Mem[ 96] = {4'h0, 4'h0, 4'h5};
        Mem[ 97] = {4'h0, 4'h0, 4'h5};
        Mem[ 98] = {4'h0, 4'h0, 4'h5};
        Mem[ 99] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[100] = {4'h0, 4'h0, 4'h5};
        Mem[101] = {4'h0, 4'h0, 4'h5};
        Mem[102] = {4'h0, 4'h0, 4'h5};
        Mem[103] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[104] = {4'h0, 4'h0, 4'h4};
        Mem[105] = {4'h0, 4'h0, 4'h4};
        Mem[106] = {4'h0, 4'h0, 4'h4};
        Mem[107] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[108] = {4'h0, 4'h0, 4'h4};
        Mem[109] = {4'h0, 4'h0, 4'h4};
        Mem[110] = {4'h0, 4'h0, 4'h4};
        Mem[111] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[112] = {4'h0, 4'h0, 4'h3};
        Mem[113] = {4'h0, 4'h0, 4'h3};
        Mem[114] = {4'h0, 4'h0, 4'h3};
        Mem[115] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[116] = {4'h0, 4'h0, 4'h3};
        Mem[117] = {4'h0, 4'h0, 4'h3};
        Mem[118] = {4'h0, 4'h0, 4'h3};
        Mem[119] = {4'h0, 4'h0, 4'h0}; // 空
        Mem[120] = {4'h0, 4'h0, 4'h2};
        Mem[121] = {4'h0, 4'h0, 4'h2};
        Mem[122] = {4'h0, 4'h0, 4'h2};
        Mem[123] = {4'h0, 4'h0, 4'h2};
        Mem[124] = {4'h0, 4'h0, 4'h2};
        Mem[125] = {4'h0, 4'h0, 4'h2};
        Mem[126] = {4'h0, 4'h0, 4'h2};
        Mem[127] = {4'h0, 4'h0, 4'h0}; // 空
    end

    assign data = Mem[addr];

endmodule